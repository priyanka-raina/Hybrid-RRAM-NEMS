.subckt cluster_0 n12849cf0 n12849cd8

m1285d4b0 n12849cf0 n12849cd8 0 0 n l=1e-07 w=1.9e-07 m=1

m1285d438 n12849cf0 n12849cd8 n12849170 n12849170 p l=1e-07 w=4.15e-07 m=1

.ends

* Finished writing spice file on Date: Mon Jun 24 06:44:47 2019

