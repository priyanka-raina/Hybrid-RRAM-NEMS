*.SCALE METER
*.LDD
.GLOBAL gnd vdd vb

***
.hdl nem_relay_4T.va

.subckt NEM4T_OFF Vsrc Vdrn
Xnem Vdrn gnd Vsrc vb Vpi=0.8 Vpo=0.2 rch=1E3 tdmec=1E-9 Cgbon=2E-17 Cgboff=1.5E-17 on_flg=0
.ends NEM4T_OFF
