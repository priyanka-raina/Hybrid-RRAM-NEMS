.title <test_4T_simple_copy0_hold.sp>

.hdl simple_rram.va
.hdl nem_relay_4T.va

** Device parameters **


** Test filamentary RRAM **
Rtfr Vlow Vhigh
Xrram_fil te be SimpleRRAM

.end